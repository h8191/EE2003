module forwarder(
	input [4:0] rs1,
	input [4:0] rs2,
	input [32:0] imm,
	input [34:0] dec_ex,
	input [34:0] ex_mem,
	input [34:0] mem_wb,

	output reg [31:0] alu_in1, alu_in2
);
	

endmodule